library verilog;
use verilog.vl_types.all;
entity mainctrl_tb is
end mainctrl_tb;
