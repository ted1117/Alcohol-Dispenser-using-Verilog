library verilog;
use verilog.vl_types.all;
entity tb_seg_top is
end tb_seg_top;
